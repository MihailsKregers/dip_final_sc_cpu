`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   22:46:52 01/20/2021
// Design Name:   computer_simulator
// Module Name:   /media/user/b70d0e4c-8ac3-4f9b-aabb-068906af6193/14.7/ISE_DS/DIP_project_processor/test_computer.v
// Project Name:  DIP_project_processor
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: computer_simulator
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module test_computer;

	// Outputs
	wire ;

	// Instantiate the Unit Under Test (UUT)
	computer_simulator uut (
		.()
	);

	initial begin
		// Initialize Inputs

		// Wait 100 ns for global reset to finish
		#100;
        
		// Add stimulus here

	end
      
endmodule

